module forwarding_unit(output	    stallF, stallD,
		       output	    forwardAD, forwardBD,
		       output	    flushE,
		       output [1:0] forwardAE, forwardBE);

endmodule
