module hazard_detector_tb;

  //[TODO:] hazard_detector testbench

endmodule
