module forwarding_unit();

//[TODO:] Ports and Implementation (Also not sure if this is designed at top level)

endmodule
