module forwwarding_unit_tb;

  //[TODO:] Forwarding Unit Testbench

endmodule
