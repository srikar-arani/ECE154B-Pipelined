module hazard_detector();

  //[TODO:] Ports and Implementation

endmodule
