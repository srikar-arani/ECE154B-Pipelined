module multiplier(input  [31:0] a,b,
		  input clk,start,is_signed,
		  output [63:0] s);

  //[TODO:] Multiplier Implementation

endmodule
